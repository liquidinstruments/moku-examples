library IEEE;
use IEEE.Std_Logic_1164.all;
use IEEE.Numeric_Std.all;


architecture Behavioural of CustomWrapper is
begin
    -- ___ <= InputA;
    -- ___ <= InputB;
    -- ___ <= InputC;
    -- ___ <= InputD;

    -- ___ <= Control(0);
    -- ___ <= Control(1);
    -- ___ <= Control(2);
    --      ...
    -- ___ <= Control(15);

    -- OutputA => ___;
    -- OutputB => ___;
    -- OutputC => ___;
    -- OutputD => ___;
    
end architecture;
